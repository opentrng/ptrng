library ieee;
use ieee.std_logic_1164.all;

package settings is
	constant T: natural := 1;
	constant RO_LEN: array (0 to T) of natural := (20, 20);
end package;
