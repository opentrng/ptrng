library ieee;
use std.textio.all;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

-- Test bench entity for COSO.
entity coso_tb is
end entity;

-- Implementation of the testbench for simulation.
architecture sim of coso_tb is

	signal ro1: std_logic := '0';
	signal ro2: std_logic := '0';

	signal coso_clk: std_logic;
	signal coso_lsb: std_logic;
	signal coso_raw: std_logic_vector (31 downto 0);

	file fout: text;

begin

	-- COSO is the design under test
	dut: entity work.coso(original)
	port map (
		ro1 => ro1,
		ro2 => ro2,
		clk => coso_clk,
		lsb => coso_lsb,
		raw => coso_raw
	);

	-- Simulation of RO1 with data generated by the RO emulator
	rofile1: entity work.rofile
	generic map (
		PATH => "../../data/ro1.txt"
	)
	port map (
		enable => '1',
		osc => ro1
	);

	-- Simulation of RO2 with data generated by the RO emulator
	rofile2: entity work.rofile
	generic map (
		PATH => "../../data/ro2.txt"
	)
	port map (
		enable => '1',
		osc => ro2
	);

	-- Write each COSO random bit to the output file 'coso.txt'
	file_open(fout, "../../data/coso_tb.txt",  write_mode);
	output: process (coso_clk)
		variable outline: line;
	begin
		if rising_edge(coso_clk) then
			write(outline, to_integer(unsigned(coso_raw)));
			writeline(fout, outline);
		end if;
	end process;

end architecture;
