library ieee;
use ieee.std_logic_1164.all;

package constants is

	-- Digitizer types
	constant TEST: natural := 0;
	constant ERO: natural := 1;
	constant MURO: natural := 2;
	constant COSO: natural := 3;

end package;
